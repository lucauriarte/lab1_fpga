-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Sat Nov 08 13:17:54 2025

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY maquina_i2c IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        SDA : IN STD_LOGIC := '0';
        fin_dir : IN STD_LOGIC := '0';
        soy : IN STD_LOGIC := '0';
        fin_dato : IN STD_LOGIC := '0';
        hab_dir : OUT STD_LOGIC;
        hab_dat : OUT STD_LOGIC;
        ack_o : OUT STD_LOGIC
    );
END maquina_i2c;

ARCHITECTURE BEHAVIOR OF maquina_i2c IS
    TYPE type_fstate IS (ocioso,Guarda_dir,R_W,ACK,Guarda_dato);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,SDA,fin_dir,soy,fin_dato)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= ocioso;
            hab_dir <= '0';
            hab_dat <= '0';
            ack_o <= '0';
        ELSE
            hab_dir <= '0';
            hab_dat <= '0';
            ack_o <= '0';
            CASE fstate IS
                WHEN ocioso =>
                    IF ((SDA = '0')) THEN
                        reg_fstate <= Guarda_dir;
                    ELSIF ((SDA = '1')) THEN
                        reg_fstate <= ocioso;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= ocioso;
                    END IF;
                WHEN Guarda_dir =>
                    IF (((fin_dir = '1') AND (soy = '0'))) THEN
                        reg_fstate <= ocioso;
                    ELSIF (((fin_dir = '1') AND (soy = '1'))) THEN
                        reg_fstate <= R_W;
                    ELSIF ((fin_dir = '0')) THEN
                        reg_fstate <= Guarda_dir;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Guarda_dir;
                    END IF;

                    hab_dir <= '1';
                WHEN R_W =>
                    reg_fstate <= ACK;
                WHEN ACK =>
                    reg_fstate <= Guarda_dato;

                    ack_o <= '1';
                WHEN Guarda_dato =>
                    IF ((fin_dato = '1')) THEN
                        reg_fstate <= ocioso;
                    ELSIF ((fin_dato = '0')) THEN
                        reg_fstate <= Guarda_dato;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Guarda_dato;
                    END IF;

                    hab_dat <= '1';
                WHEN OTHERS => 
                    hab_dir <= 'X';
                    hab_dat <= 'X';
                    ack_o <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
