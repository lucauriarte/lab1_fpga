-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition"
-- CREATED		"Thu Nov 06 16:39:54 2025"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY parte_c IS 
	PORT
	(
		A0 :  IN  STD_LOGIC;
		B0 :  IN  STD_LOGIC;
		A1 :  IN  STD_LOGIC;
		B1 :  IN  STD_LOGIC;
		CLK :  IN  STD_LOGIC;
		P0 :  OUT  STD_LOGIC;
		P1 :  OUT  STD_LOGIC;
		P2 :  OUT  STD_LOGIC;
		P3 :  OUT  STD_LOGIC;
		Signo :  OUT  STD_LOGIC;
		Cero :  OUT  STD_LOGIC
	);
END parte_c;

ARCHITECTURE bdf_type OF parte_c IS 

COMPONENT parte_a
	PORT(A : IN STD_LOGIC;
		 B : IN STD_LOGIC;
		 Cin : IN STD_LOGIC;
		 S : OUT STD_LOGIC;
		 Cout : OUT STD_LOGIC
	);
END COMPONENT;

SIGNAL	C0 :  STD_LOGIC;
SIGNAL	C1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_24 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_25 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_26 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_27 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_28 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_29 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_30 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_31 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_32 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_33 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC;


BEGIN 
SYNTHESIZED_WIRE_4 <= '1';
SYNTHESIZED_WIRE_6 <= '0';
SYNTHESIZED_WIRE_19 <= '0';




PROCESS(CLK)
BEGIN
IF (RISING_EDGE(CLK)) THEN
	SYNTHESIZED_WIRE_26 <= A0;
END IF;
END PROCESS;


b2v_inst11 : parte_a
PORT MAP(A => SYNTHESIZED_WIRE_24,
		 B => SYNTHESIZED_WIRE_1,
		 Cin => SYNTHESIZED_WIRE_2,
		 S => SYNTHESIZED_WIRE_31);


PROCESS(CLK)
BEGIN
IF (RISING_EDGE(CLK)) THEN
	SYNTHESIZED_WIRE_32 <= B0;
END IF;
END PROCESS;


PROCESS(CLK)
BEGIN
IF (RISING_EDGE(CLK)) THEN
	SYNTHESIZED_WIRE_28 <= A1;
END IF;
END PROCESS;


PROCESS(CLK)
BEGIN
IF (RISING_EDGE(CLK)) THEN
	SYNTHESIZED_WIRE_33 <= B1;
END IF;
END PROCESS;


PROCESS(CLK)
BEGIN
IF (RISING_EDGE(CLK)) THEN
	P0 <= SYNTHESIZED_WIRE_25;
END IF;
END PROCESS;


b2v_inst16 : parte_a
PORT MAP(A => SYNTHESIZED_WIRE_4,
		 B => SYNTHESIZED_WIRE_5,
		 Cin => SYNTHESIZED_WIRE_6,
		 S => C0);



SYNTHESIZED_WIRE_5 <= NOT(SYNTHESIZED_WIRE_26);




b2v_inst20 : parte_a
PORT MAP(A => C0,
		 B => SYNTHESIZED_WIRE_27,
		 S => C1);


SYNTHESIZED_WIRE_27 <= NOT(SYNTHESIZED_WIRE_28);



PROCESS(CLK)
BEGIN
IF (RISING_EDGE(CLK)) THEN
	P1 <= SYNTHESIZED_WIRE_29;
END IF;
END PROCESS;


PROCESS(CLK)
BEGIN
IF (RISING_EDGE(CLK)) THEN
	P2 <= SYNTHESIZED_WIRE_30;
END IF;
END PROCESS;


PROCESS(CLK)
BEGIN
IF (RISING_EDGE(CLK)) THEN
	P3 <= SYNTHESIZED_WIRE_31;
END IF;
END PROCESS;


PROCESS(CLK)
BEGIN
IF (RISING_EDGE(CLK)) THEN
	Signo <= SYNTHESIZED_WIRE_31;
END IF;
END PROCESS;


SYNTHESIZED_WIRE_16 <= NOT(SYNTHESIZED_WIRE_31 OR SYNTHESIZED_WIRE_29 OR SYNTHESIZED_WIRE_30 OR SYNTHESIZED_WIRE_25);


PROCESS(CLK)
BEGIN
IF (RISING_EDGE(CLK)) THEN
	Cero <= SYNTHESIZED_WIRE_16;
END IF;
END PROCESS;


b2v_inst3 : parte_a
PORT MAP(A => SYNTHESIZED_WIRE_17,
		 B => SYNTHESIZED_WIRE_24,
		 Cin => SYNTHESIZED_WIRE_19,
		 S => SYNTHESIZED_WIRE_29,
		 Cout => SYNTHESIZED_WIRE_22);


SYNTHESIZED_WIRE_25 <= SYNTHESIZED_WIRE_26 AND SYNTHESIZED_WIRE_32;


SYNTHESIZED_WIRE_24 <= SYNTHESIZED_WIRE_28 AND SYNTHESIZED_WIRE_32;


SYNTHESIZED_WIRE_17 <= C0 AND SYNTHESIZED_WIRE_33;


b2v_inst7 : parte_a
PORT MAP(A => SYNTHESIZED_WIRE_24,
		 B => SYNTHESIZED_WIRE_21,
		 Cin => SYNTHESIZED_WIRE_22,
		 S => SYNTHESIZED_WIRE_30,
		 Cout => SYNTHESIZED_WIRE_2);


SYNTHESIZED_WIRE_21 <= SYNTHESIZED_WIRE_33 AND C1;


SYNTHESIZED_WIRE_1 <= SYNTHESIZED_WIRE_33 AND SYNTHESIZED_WIRE_27;


END bdf_type;