-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Fri Nov 07 14:15:39 2025

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY parte_e IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        x : IN STD_LOGIC := '0';
        z : OUT STD_LOGIC_VECTOR(0 TO 3)
    );
END parte_e;

ARCHITECTURE BEHAVIOR OF parte_e IS
    TYPE type_fstate IS (state1,state2,state3,state4,state5,state6,state7,state8);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,x)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= state1;
            z <= "0000";
        ELSE
            z <= "0000";
            CASE fstate IS
                WHEN state1 =>
                    IF ((x = '0')) THEN
                        reg_fstate <= state2;
                    ELSIF ((x = '1')) THEN
                        reg_fstate <= state5;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state1;
                    END IF;

                    z <= "0000";
                WHEN state2 =>
                    reg_fstate <= state3;

                    z <= "0110";
                WHEN state3 =>
                    IF ((x = '0')) THEN
                        reg_fstate <= state4;
                    ELSIF ((x = '1')) THEN
                        reg_fstate <= state7;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state3;
                    END IF;

                    z <= "1111";
                WHEN state4 =>
                    reg_fstate <= state8;

                    z <= "1001";
                WHEN state5 =>
                    reg_fstate <= state6;

                    z <= "1000";
                WHEN state6 =>
                    reg_fstate <= state3;

                    z <= "1100";
                WHEN state7 =>
                    reg_fstate <= state8;

                    z <= "1110";
                WHEN state8 =>
                    reg_fstate <= state1;

                    z <= "0000";
                WHEN OTHERS => 
                    z <= "XXXX";
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
